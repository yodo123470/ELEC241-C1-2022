module task3;

//Write solution here

endmodule
