module task3_tb;

//Write testbench here

endmodule
